`timescale 1ns / 1ns
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 24.05.2022 19:18:39
// Design Name: 
// Module Name: censor_rtl_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module censor_rtl_tb();
    
    int i = 0;
    
    reg clock, reset, bloom_write, data_ready, enable;
    reg string_end = 0;
    reg [7:0] char_in;
    reg [7:0] char_out;
    reg [0:1016][7:0] tab_char_in = {   8'h41, 8'h67, 8'h65, 8'h6e, 8'h74, 8'h73, 8'h20, 8'h73, 8'h65, 8'h72, 8'h69, 8'h65, 8'h73, 8'h20, 8'h54, 8'h75, 8'h67, 8'h6f,
                                        8'h72, 8'h20, 8'h61, 8'h67, 8'h65, 8'h6e, 8'h74, 8'h20, 8'h54, 8'h68, 8'h65, 8'h20, 8'h50, 8'h68, 8'h61, 8'h6e, 8'h74, 8'h6f,
                                        8'h6d, 8'h20, 8'h41, 8'h67, 8'h65, 8'h6e, 8'h74, 8'h73, 8'h20, 8'h77, 8'h65, 8'h72, 8'h65, 8'h20, 8'h61, 8'h72, 8'h6d, 8'h65, 
                                        8'h64, 8'h20, 8'h77, 8'h69, 8'h74, 8'h68, 8'h20, 8'h6e, 8'h69, 8'h6e, 8'h6a, 8'h61, 8'h20, 8'h77, 8'h65, 8'h61, 8'h70, 8'h6f, 
                                        8'h6e, 8'h73, 8'h20, 8'h73, 8'h75, 8'h63, 8'h68, 8'h20, 8'h61, 8'h73, 8'h20, 8'h73, 8'h68, 8'h75, 8'h72, 8'h69, 8'h6b, 8'h65, 
                                        8'h6e, 8'h20, 8'h61, 8'h6e, 8'h64, 8'h20, 8'h75, 8'h73, 8'h65, 8'h64, 8'h20, 8'h67, 8'h75, 8'h6e, 8'h73, 8'h20, 8'h22, 8'h6f, 
                                        8'h6e, 8'h6c, 8'h79, 8'h20, 8'h61, 8'h73, 8'h20, 8'h61, 8'h20, 8'h6c, 8'h61, 8'h73, 8'h74, 8'h20, 8'h72, 8'h65, 8'h73, 8'h6f, 
                                        8'h72, 8'h74, 8'h2c, 8'h22, 8'h20, 8'h61, 8'h73, 8'h20, 8'h77, 8'h61, 8'h73, 8'h20, 8'h70, 8'h61, 8'h74, 8'h69, 8'h65, 8'h6e, 
                                        8'h74, 8'h6c, 8'h79, 8'h20, 8'h65, 8'h78, 8'h70, 8'h6c, 8'h61, 8'h69, 8'h6e, 8'h65, 8'h64, 8'h20, 8'h74, 8'h6f, 8'h20, 8'h74, 
                                        8'h68, 8'h65, 8'h20, 8'h6f, 8'h6e, 8'h6c, 8'h79, 8'h20, 8'h66, 8'h65, 8'h6d, 8'h61, 8'h6c, 8'h65, 8'h20, 8'h6d, 8'h65, 8'h6d, 
                                        8'h62, 8'h65, 8'h72, 8'h20, 8'h69, 8'h6e, 8'h20, 8'h74, 8'h68, 8'h65, 8'h20, 8'h74, 8'h69, 8'h74, 8'h6c, 8'h65, 8'h20, 8'h73, 
                                        8'h65, 8'h71, 8'h75, 8'h65, 8'h6e, 8'h63, 8'h65, 8'h20, 8'h6f, 8'h66, 8'h20, 8'h65, 8'h61, 8'h63, 8'h68, 8'h20, 8'h65, 8'h70, 
                                        8'h69, 8'h73, 8'h6f, 8'h64, 8'h65, 8'h2e, 8'h20, 8'h54, 8'h68, 8'h65, 8'h79, 8'h20, 8'h68, 8'h61, 8'h64, 8'h20, 8'h74, 8'h68, 
                                        8'h65, 8'h20, 8'h61, 8'h62, 8'h69, 8'h6c, 8'h69, 8'h74, 8'h79, 8'h20, 8'h74, 8'h6f, 8'h20, 8'h6a, 8'h75, 8'h6d, 8'h70, 8'h20, 
                                        8'h62, 8'h61, 8'h63, 8'h6b, 8'h77, 8'h61, 8'h72, 8'h64, 8'h73, 8'h20, 8'h75, 8'h70, 8'h20, 8'h6f, 8'h6e, 8'h74, 8'h6f, 8'h20, 
                                        8'h74, 8'h68, 8'h65, 8'h20, 8'h6c, 8'h69, 8'h6d, 8'h62, 8'h73, 8'h20, 8'h6f, 8'h66, 8'h20, 8'h74, 8'h72, 8'h65, 8'h65, 8'h73, 
                                        8'h20, 8'h61, 8'h6e, 8'h64, 8'h20, 8'h63, 8'h6f, 8'h75, 8'h6c, 8'h64, 8'h20, 8'h68, 8'h6f, 8'h6c, 8'h64, 8'h20, 8'h61, 8'h20, 
                                        8'h70, 8'h69, 8'h65, 8'h63, 8'h65, 8'h20, 8'h6f, 8'h66, 8'h20, 8'h63, 8'h6c, 8'h6f, 8'h74, 8'h68, 8'h20, 8'h77, 8'h69, 8'h74, 
                                        8'h68, 8'h20, 8'h61, 8'h20, 8'h62, 8'h72, 8'h69, 8'h63, 8'h6b, 8'h20, 8'h70, 8'h61, 8'h74, 8'h74, 8'h65, 8'h72, 8'h6e, 8'h20, 
                                        8'h6f, 8'h6e, 8'h20, 8'h69, 8'h74, 8'h20, 8'h69, 8'h6e, 8'h20, 8'h66, 8'h72, 8'h6f, 8'h6e, 8'h74, 8'h20, 8'h6f, 8'h66, 8'h20, 
                                        8'h74, 8'h68, 8'h65, 8'h6d, 8'h20, 8'h61, 8'h6e, 8'h64, 8'h20, 8'h74, 8'h68, 8'h75, 8'h73, 8'h20, 8'h62, 8'h6c, 8'h65, 8'h6e, 
                                        8'h64, 8'h20, 8'h69, 8'h6e, 8'h74, 8'h6f, 8'h20, 8'h74, 8'h68, 8'h65, 8'h20, 8'h77, 8'h61, 8'h6c, 8'h6c, 8'h20, 8'h62, 8'h65, 
                                        8'h68, 8'h69, 8'h6e, 8'h64, 8'h20, 8'h74, 8'h68, 8'h65, 8'h6d, 8'h2c, 8'h20, 8'h62, 8'h65, 8'h63, 8'h6f, 8'h6d, 8'h69, 8'h6e, 
                                        8'h67, 8'h20, 8'h69, 8'h6e, 8'h76, 8'h69, 8'h73, 8'h69, 8'h62, 8'h6c, 8'h65, 8'h20, 8'h74, 8'h6f, 8'h20, 8'h74, 8'h68, 8'h65, 
                                        8'h69, 8'h72, 8'h20, 8'h6f, 8'h70, 8'h70, 8'h6f, 8'h6e, 8'h65, 8'h6e, 8'h74, 8'h73, 8'h2e, 8'h20, 8'h54, 8'h68, 8'h65, 8'h20, 
                                        8'h73, 8'h65, 8'h72, 8'h69, 8'h65, 8'h73, 8'h20, 8'h73, 8'h74, 8'h61, 8'h72, 8'h72, 8'h65, 8'h64, 8'h20, 8'h4a, 8'h6f, 8'h68, 
                                        8'h20, 8'h4d, 8'h69, 8'h7a, 8'h75, 8'h6b, 8'h69, 8'h20, 8'h61, 8'h73, 8'h20, 8'h50, 8'h68, 8'h61, 8'h6e, 8'h74, 8'h61, 8'h72, 
                                        8'h2c, 8'h20, 8'h74, 8'h68, 8'h65, 8'h20, 8'h6c, 8'h65, 8'h61, 8'h64, 8'h65, 8'h72, 8'h20, 8'h6f, 8'h66, 8'h20, 8'h74, 8'h68, 
                                        8'h65, 8'h20, 8'h50, 8'h68, 8'h61, 8'h6e, 8'h74, 8'h6f, 8'h6d, 8'h20, 8'h41, 8'h67, 8'h65, 8'h6e, 8'h74, 8'h73, 8'h20, 8'h4f, 
                                        8'h74, 8'h68, 8'h65, 8'h72, 8'h20, 8'h41, 8'h67, 8'h65, 8'h6e, 8'h74, 8'h73, 8'h20, 8'h69, 8'h6e, 8'h63, 8'h6c, 8'h75, 8'h64, 
                                        8'h65, 8'h64, 8'h20, 8'h54, 8'h75, 8'h67, 8'h6f, 8'h72, 8'h20, 8'h43, 8'h6f, 8'h72, 8'h64, 8'h6f, 8'h2c, 8'h20, 8'h5a, 8'h65, 
                                        8'h6d, 8'h6f, 8'h20, 8'h61, 8'h6e, 8'h64, 8'h20, 8'h61, 8'h20, 8'h66, 8'h65, 8'h6d, 8'h61, 8'h6c, 8'h65, 8'h20, 8'h61, 8'h67, 
                                        8'h65, 8'h6e, 8'h74, 8'h20, 8'h2c, 8'h20, 8'h4d, 8'h61, 8'h72, 8'h67, 8'h6f, 8'h20, 8'h28, 8'h6c, 8'h61, 8'h74, 8'h65, 8'h72, 
                                        8'h20, 8'h72, 8'h65, 8'h70, 8'h6c, 8'h61, 8'h63, 8'h65, 8'h64, 8'h20, 8'h62, 8'h79, 8'h20, 8'h47, 8'h69, 8'h6e, 8'h61, 8'h29, 
                                        8'h2e, 8'h20, 8'h54, 8'h68, 8'h65, 8'h72, 8'h65, 8'h20, 8'h77, 8'h61, 8'h73, 8'h20, 8'h61, 8'h6c, 8'h73, 8'h6f, 8'h20, 8'h61, 
                                        8'h20, 8'h73, 8'h6d, 8'h61, 8'h6c, 8'h6c, 8'h20, 8'h62, 8'h6f, 8'h79, 8'h20, 8'h61, 8'h67, 8'h65, 8'h6e, 8'h74, 8'h20, 8'h2c, 
                                        8'h20, 8'h54, 8'h6f, 8'h6d, 8'h62, 8'h61, 8'h20, 8'h4f, 8'h74, 8'h68, 8'h65, 8'h72, 8'h20, 8'h41, 8'h67, 8'h65, 8'h6e, 8'h74, 
                                        8'h73, 8'h20, 8'h74, 8'h68, 8'h61, 8'h74, 8'h20, 8'h6a, 8'h6f, 8'h69, 8'h6e, 8'h65, 8'h64, 8'h20, 8'h6c, 8'h61, 8'h74, 8'h65, 
                                        8'h72, 8'h20, 8'h69, 8'h6e, 8'h20, 8'h74, 8'h68, 8'h65, 8'h20, 8'h73, 8'h65, 8'h72, 8'h69, 8'h65, 8'h73, 8'h20, 8'h77, 8'h65, 
                                        8'h72, 8'h65, 8'h20, 8'h41, 8'h6e, 8'h64, 8'h61, 8'h72, 8'h20, 8'h28, 8'h77, 8'h68, 8'h6f, 8'h20, 8'h73, 8'h65, 8'h65, 8'h6d, 
                                        8'h65, 8'h64, 8'h20, 8'h74, 8'h6f, 8'h20, 8'h72, 8'h65, 8'h70, 8'h6c, 8'h61, 8'h63, 8'h65, 8'h20, 8'h54, 8'h75, 8'h67, 8'h6f, 
                                        8'h72, 8'h20, 8'h29, 8'h20, 8'h61, 8'h6e, 8'h64, 8'h20, 8'h4d, 8'h75, 8'h6e, 8'h64, 8'h6f, 8'h2c, 8'h20, 8'h77, 8'h68, 8'h6f, 
                                        8'h20, 8'h63, 8'h6f, 8'h75, 8'h6c, 8'h64, 8'h20, 8'h72, 8'h6f, 8'h6c, 8'h6c, 8'h20, 8'h68, 8'h69, 8'h6d, 8'h73, 8'h65, 8'h6c, 
                                        8'h66, 8'h20, 8'h75, 8'h70, 8'h20, 8'h69, 8'h6e, 8'h74, 8'h6f, 8'h20, 8'h61, 8'h20, 8'h62, 8'h6f, 8'h77, 8'h6c, 8'h69, 8'h6e, 
                                        8'h67, 8'h20, 8'h62, 8'h61, 8'h6c, 8'h6c, 8'h20, 8'h74, 8'h6f, 8'h20, 8'h6b, 8'h6e, 8'h6f, 8'h63, 8'h6b, 8'h20, 8'h6f, 8'h76, 
                                        8'h65, 8'h72, 8'h20, 8'h74, 8'h68, 8'h65, 8'h20, 8'h76, 8'h69, 8'h6c, 8'h6c, 8'h61, 8'h69, 8'h6e, 8'h73, 8'h2e, 8'h20, 8'h54, 
                                        8'h75, 8'h67, 8'h6f, 8'h72, 8'h20, 8'h77, 8'h61, 8'h73, 8'h20, 8'h6b, 8'h69, 8'h6c, 8'h6c, 8'h65, 8'h64, 8'h20, 8'h62, 8'h79, 
                                        8'h20, 8'h61, 8'h20, 8'h62, 8'h6f, 8'h6d, 8'h62, 8'h20, 8'h69, 8'h6e, 8'h20, 8'h6f, 8'h6e, 8'h65, 8'h20, 8'h6f, 8'h66, 8'h20, 
                                        8'h74, 8'h68, 8'h65, 8'h20, 8'h65, 8'h70, 8'h69, 8'h73, 8'h6f, 8'h64, 8'h65, 8'h73, 8'h2c, 8'h20, 8'h6c, 8'h65, 8'h61, 8'h76, 
                                        8'h69, 8'h6e, 8'h67, 8'h20, 8'h62, 8'h65, 8'h68, 8'h69, 8'h6e, 8'h64, 8'h20, 8'h6f, 8'h6e, 8'h6c, 8'h79, 8'h20, 8'h61, 8'h20, 
                                        8'h62, 8'h6f, 8'h6f, 8'h74, 8'h20, 8'h74, 8'h68, 8'h61, 8'h74, 8'h20, 8'h6d, 8'h61, 8'h6e, 8'h79, 8'h20, 8'h66, 8'h61, 8'h6e, 
                                        8'h73, 8'h20, 8'h72, 8'h65, 8'h6d, 8'h65, 8'h6d, 8'h62, 8'h65, 8'h72, 8'h20, 8'h61, 8'h73, 8'h20, 8'h61, 8'h20, 8'h73, 8'h61, 
                                        8'h64, 8'h20, 8'h6d, 8'h6f, 8'h6d, 8'h65, 8'h6e, 8'h74, 8'h20, 8'h69, 8'h6e, 8'h20, 8'h74, 8'h68, 8'h65, 8'h20, 8'h73, 8'h65, 
                                        8'h72, 8'h69, 8'h65, 8'h73, 8'h20, 8'h2e, 8'h20, 8'h41, 8'h6e, 8'h6f, 8'h74, 8'h68, 8'h65, 8'h72, 8'h20, 8'h61, 8'h67, 8'h65, 
                                        8'h6e, 8'h74, 8'h20, 8'h2c, 8'h20, 8'h47, 8'h69, 8'h6e, 8'h6f, 8'h2c, 8'h20, 8'h77, 8'h61, 8'h73, 8'h20, 8'h6b, 8'h69, 8'h6c, 
                                        8'h6c, 8'h65, 8'h64, 8'h20, 8'h69, 8'h6e, 8'h20, 8'h74, 8'h68, 8'h65, 8'h20, 8'h66, 8'h69, 8'h72, 8'h73, 8'h74, 8'h20, 8'h65, 
                                        8'h70, 8'h69, 8'h73, 8'h6f, 8'h64, 8'h65, 8'h2e, 8'h20 };
    
    censor_rtl censor(clock, reset, enable, bloom_write, char_in, char_out, data_ready);

    //Clock generator
    initial
     clock <= 1'b0;
    always
     #50 clock <= ~clock;
    
    //Reset signal
    initial
    begin
     reset <= 1'b1;
     #100 reset <= 1'b0;
    end
    
    //enable signal
    initial
    begin
        enable <= 1'b1;
        #9700 enable <= 1'b0;
        #1000 enable <= 1'b1;
    end
    
    //write signal
    initial
    begin
     bloom_write <= 1'b1;
     #2700 bloom_write <= 1'b0;
    end
    
    //Data in
    always @ (negedge clock) begin
        char_in = tab_char_in[i];
        i++;
        i = i%1017;
        if(i == 1016)
            string_end <= ~string_end;       
    end

endmodule
